module id_ex

import rv32i_types::*;
(
    input clk,
    input rst,


    input rv32i_word pc_reg_in,
    input rv32i_word reg_1_in,
    input rv32i_word reg_2_in,
    input rv32i_reg reg_dest_in,
    input rv32i_control_word cntrl_word_in,
    input logic [2:0] funct3_in,
    input stall,
	input flush,
    input rv32i_word i_imm_in,
    input rv32i_word s_imm_in,
    input rv32i_word b_imm_in,
    input rv32i_word u_imm_in,
    input rv32i_word j_imm_in,
    input logic stall_nop,
    input rv32i_reg rs1_id_in,
    input rv32i_reg rs2_id_in,
	input logic br_pred_in,
	output logic br_pred_out,
	input rv32i_word br_pred_pc_in,
	output rv32i_word br_pred_pc_out,

    output rv32i_word i_imm_out,
    output rv32i_word s_imm_out,
    output rv32i_word b_imm_out,
    output rv32i_word u_imm_out,
    output rv32i_word j_imm_out,
    output rv32i_control_word cntrl_word_out,
    output logic [2:0] funct3_out,
    output rv32i_reg reg_dest_out,
    output rv32i_word reg_1_out,
    output rv32i_word reg_2_out,
    output rv32i_word pc_reg_out,
    output rv32i_reg rs1_id_out,
    output rv32i_reg rs2_id_out,


	input rv32i_opcode opcode_in,
	output rv32i_opcode opcode_out
);

//assign opcode_out = opcode_in;

always_ff @(posedge clk) begin
    if (rst) begin
        pc_reg_out <= rv32i_word'(32'b0);
        reg_1_out <= rv32i_word'(32'b0);
        reg_2_out <=rv32i_word'(32'b0);
        reg_dest_out <= rv32i_reg'(5'b0); //may need to change later cuase this is "reg0"
        i_imm_out <= rv32i_word'(32'b0);
        s_imm_out <= rv32i_word'(32'b0);
        b_imm_out <= rv32i_word'(32'b0);
        u_imm_out <= rv32i_word'(32'b0);
        j_imm_out <= rv32i_word'(32'b0);
        cntrl_word_out <= rv32i_control_word'(1'b0); //fix when size of control word is known
        funct3_out <= 3'b0;
		opcode_out <= opcode_in;
        rs1_id_out <= rv32i_reg'(1'b0);
        rs2_id_out <= rv32i_reg'(1'b0);
		br_pred_out <= 1'b0;
		br_pred_pc_out <= rv32i_word'(32'b0);
    end
	else if (flush /*|| (flush && stall_nop) || (flush && stall)*/) begin
		//opcode_out <= rv32i_opcode'(7'h13); //if not stalling replace no-op to prevent double branch.
		//cntrl_word_out <= rv32i_control_word'(1'b0);
            cntrl_word_out <= rv32i_control_word'({3'b0,3'b0,1'b0,2'b0, 3'b0, 4'b0, 2'b0, 1'b0, 1'b0, 1'b1, 7'h13});
            pc_reg_out <= rv32i_word'(32'b0);
            reg_1_out <= rv32i_word'(32'b0);
            reg_2_out <=rv32i_word'(32'b0);
            reg_dest_out <= rv32i_reg'(5'b0); //may need to change later cuase this is "reg0"
            i_imm_out <= rv32i_word'(32'b0);
            s_imm_out <= rv32i_word'(32'b0);
            b_imm_out <= rv32i_word'(32'b0);
            u_imm_out <= rv32i_word'(32'b0);
            j_imm_out <= rv32i_word'(32'b0);
            cntrl_word_out <= rv32i_control_word'(1'b0); //fix when size of control word is known
            funct3_out <= 3'b0;
		    opcode_out <= rv32i_opcode'(7'h13);
            rs1_id_out <= rv32i_reg'(1'b0);
            rs2_id_out <= rv32i_reg'(1'b0);
	end
    else begin
        if (~stall) begin
            pc_reg_out <=pc_reg_in; 
            reg_1_out <= reg_1_in;
            reg_2_out <=reg_2_in;
            reg_dest_out <= reg_dest_in;
            i_imm_out <= i_imm_in;
            s_imm_out <= s_imm_in;
            b_imm_out <= b_imm_in;
            u_imm_out <= u_imm_in;
            j_imm_out <= j_imm_in;
            cntrl_word_out <= cntrl_word_in;
            funct3_out <= funct3_in; 
		    opcode_out <= opcode_in;
            rs1_id_out <= rs1_id_in;
            rs2_id_out <= rs2_id_in;
			br_pred_out <= br_pred_in;
		   	br_pred_pc_out <= br_pred_pc_in;	
        end
        if (stall_nop) begin
            //  cntrl_word_out <= rv32i_control_word'(1'b0); //fix when size of control word is known
            cntrl_word_out <= rv32i_control_word'({3'b0,3'b0,1'b0,2'b0, 3'b0, 4'b0, 2'b0, 1'b0, 1'b0, 1'b1, 7'h13});
            pc_reg_out <= rv32i_word'(32'b0);
            reg_1_out <= rv32i_word'(32'b0);
            reg_2_out <=rv32i_word'(32'b0);
            reg_dest_out <= rv32i_reg'(5'b0); //may need to change later cuase this is "reg0"
            i_imm_out <= rv32i_word'(32'b0);
            s_imm_out <= rv32i_word'(32'b0);
            b_imm_out <= rv32i_word'(32'b0);
            u_imm_out <= rv32i_word'(32'b0);
            j_imm_out <= rv32i_word'(32'b0);
            //cntrl_word_out <= rv32i_control_word'(1'b0); //fix when size of control word is known
            funct3_out <= 3'b0;
		    opcode_out <= rv32i_opcode'(7'h13);
            rs1_id_out <= rv32i_reg'(1'b0);
            rs2_id_out <= rv32i_reg'(1'b0);
			br_pred_out <= 1'b0;
			br_pred_pc_out <= rv32i_word'(32'b0);
        end 
    end

end
endmodule : id_ex
