/************************************

	PLEASE IGNORE THIS FILE RIGHT NOW. NOT USING THIS AT ALL

*************************************/
module cpu_datapath

import rv32i_types::*;
(
	// inputs from 
	
	
	// outputs from 
);

/******** STAGE AND PIPELINE REG MODULES ********/









/******** MUXES ********/



endmodule : cpu_datapath
